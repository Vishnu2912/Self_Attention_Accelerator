package Tb;

import Acc::*;

(*synthesize*)
module mkTb(Empty);

    Ifc_load_inp dut <- mkAcc;
    Reg#(Int#(4)) start1 <- mkReg(0);   //counters
    Reg#(Int#(7)) stepq <- mkReg(0);
    Reg#(Int#(7)) stepx <- mkReg(0);

    //Parameters
    Integer in_rows = 4;
    Integer in_cols = 64;
    Integer w_cols = 16;

    //Declaration of Matrices
    Int#(64) x[in_rows][in_cols];
    Int#(64) wq[in_cols][w_cols];
    Int#(64) wk[in_cols][w_cols];
    Int#(64) wv[in_cols][w_cols];
    
    //Initialization of the Input and Weight Matrices with Quantized Integers
    
    x[0][0] = -14; x[0][1] = 11; x[0][2] = 14; x[0][3] = -16; x[0][4] = -3; x[0][5] = 13; x[0][6] = 15; x[0][7] = 1; x[0][8] = -6; x[0][9] = -14; x[0][10] = 15; x[0][11] = 4; x[0][12] = -12; x[0][13] = -1; x[0][14] = 7; x[0][15] = -14; x[0][16] = 10; x[0][17] = -8; x[0][18] = 6; x[0][19] = 8; x[0][20] = 10; x[0][21] = 2; x[0][22] = 0; x[0][23] = 13; x[0][24] = -5; x[0][25] = 3; x[0][26] = 7; x[0][27] = -8; x[0][28] = 13; x[0][29] = -1; x[0][30] = 12; x[0][31] = 8; x[0][32] = -14; x[0][33] = -16; x[0][34] = -1; x[0][35] = -8; x[0][36] = -4; x[0][37] = 3; x[0][38] = 7; x[0][39] = -1; x[0][40] = 4; x[0][41] = 12; x[0][42] = 11; x[0][43] = 14; x[0][44] = -12; x[0][45] = 4; x[0][46] = 16; x[0][47] = -6; x[0][48] = -2; x[0][49] = 10; x[0][50] = -1; x[0][51] = -14; x[0][52] = -14; x[0][53] = 15; x[0][54] = 3; x[0][55] = -12; x[0][56] = -11; x[0][57] = -7; x[0][58] = 8; x[0][59] = 7; x[0][60] = -7; x[0][61] = -9; x[0][62] = -10; x[0][63] = 12; 
x[1][0] = -6; x[1][1] = -4; x[1][2] = 6; x[1][3] = 11; x[1][4] = 10; x[1][5] = 12; x[1][6] = -1; x[1][7] = 1; x[1][8] = -7; x[1][9] = -5; x[1][10] = -9; x[1][11] = 1; x[1][12] = 13; x[1][13] = 3; x[1][14] = -6; x[1][15] = -5; x[1][16] = -5; x[1][17] = 14; x[1][18] = 6; x[1][19] = 4; x[1][20] = 11; x[1][21] = -2; x[1][22] = -16; x[1][23] = -14; x[1][24] = 5; x[1][25] = 4; x[1][26] = -1; x[1][27] = -11; x[1][28] = 0; x[1][29] = 12; x[1][30] = 9; x[1][31] = -6; x[1][32] = 8; x[1][33] = 15; x[1][34] = -1; x[1][35] = 1; x[1][36] = 14; x[1][37] = 15; x[1][38] = -12; x[1][39] = -6; x[1][40] = 15; x[1][41] = 13; x[1][42] = 9; x[1][43] = -8; x[1][44] = 10; x[1][45] = 6; x[1][46] = 8; x[1][47] = 15; x[1][48] = -6; x[1][49] = 12; x[1][50] = -10; x[1][51] = 10; x[1][52] = -14; x[1][53] = -16; x[1][54] = 12; x[1][55] = -12; x[1][56] = -13; x[1][57] = 6; x[1][58] = -11; x[1][59] = -7; x[1][60] = -10; x[1][61] = 13; x[1][62] = 15; x[1][63] = -8; 
x[2][0] = 13; x[2][1] = 11; x[2][2] = 16; x[2][3] = 12; x[2][4] = 5; x[2][5] = 0; x[2][6] = 13; x[2][7] = 11; x[2][8] = 5; x[2][9] = -7; x[2][10] = -1; x[2][11] = 4; x[2][12] = -14; x[2][13] = -4; x[2][14] = 14; x[2][15] = -15; x[2][16] = -9; x[2][17] = 2; x[2][18] = 11; x[2][19] = -1; x[2][20] = 2; x[2][21] = -11; x[2][22] = -14; x[2][23] = -10; x[2][24] = 2; x[2][25] = -6; x[2][26] = 14; x[2][27] = -7; x[2][28] = 7; x[2][29] = 9; x[2][30] = -4; x[2][31] = 6; x[2][32] = -5; x[2][33] = -11; x[2][34] = -4; x[2][35] = 11; x[2][36] = -3; x[2][37] = -10; x[2][38] = 3; x[2][39] = 13; x[2][40] = 11; x[2][41] = 12; x[2][42] = -3; x[2][43] = 1; x[2][44] = 7; x[2][45] = -9; x[2][46] = -16; x[2][47] = -3; x[2][48] = 11; x[2][49] = 10; x[2][50] = 8; x[2][51] = -4; x[2][52] = -12; x[2][53] = 11; x[2][54] = -11; x[2][55] = -13; x[2][56] = 6; x[2][57] = 0; x[2][58] = 7; x[2][59] = 13; x[2][60] = 11; x[2][61] = -4; x[2][62] = 2; x[2][63] = 13; 
x[3][0] = 2; x[3][1] = 16; x[3][2] = 15; x[3][3] = 16; x[3][4] = 0; x[3][5] = 9; x[3][6] = 12; x[3][7] = 5; x[3][8] = 6; x[3][9] = 1; x[3][10] = 14; x[3][11] = 12; x[3][12] = 14; x[3][13] = 14; x[3][14] = -11; x[3][15] = 7; x[3][16] = 9; x[3][17] = -6; x[3][18] = 10; x[3][19] = -12; x[3][20] = 3; x[3][21] = -15; x[3][22] = 4; x[3][23] = 4; x[3][24] = -12; x[3][25] = 9; x[3][26] = 7; x[3][27] = 2; x[3][28] = -5; x[3][29] = -1; x[3][30] = -6; x[3][31] = 3; x[3][32] = -10; x[3][33] = -13; x[3][34] = -2; x[3][35] = -12; x[3][36] = 10; x[3][37] = -4; x[3][38] = 12; x[3][39] = -15; x[3][40] = 9; x[3][41] = -4; x[3][42] = 5; x[3][43] = -4; x[3][44] = 4; x[3][45] = -13; x[3][46] = -13; x[3][47] = -14; x[3][48] = 7; x[3][49] = 9; x[3][50] = 4; x[3][51] = -6; x[3][52] = -6; x[3][53] = -9; x[3][54] = 6; x[3][55] = -6; x[3][56] = -15; x[3][57] = 16; x[3][58] = 6; x[3][59] = -11; x[3][60] = 9; x[3][61] = 12; x[3][62] = 6; x[3][63] = -13; 

wq[0][0] = -7; wq[0][1] = 12; wq[0][2] = 6; wq[0][3] = 16; wq[0][4] = -4; wq[0][5] = -7; wq[0][6] = -4; wq[0][7] = 8; wq[0][8] = -6; wq[0][9] = -13; wq[0][10] = 7; wq[0][11] = -14; wq[0][12] = -12; wq[0][13] = 15; wq[0][14] = 9; wq[0][15] = -14; 
wq[1][0] = 10; wq[1][1] = 9; wq[1][2] = -9; wq[1][3] = 11; wq[1][4] = -10; wq[1][5] = -1; wq[1][6] = -6; wq[1][7] = -10; wq[1][8] = -10; wq[1][9] = 2; wq[1][10] = -4; wq[1][11] = 9; wq[1][12] = 11; wq[1][13] = -13; wq[1][14] = 14; wq[1][15] = -3; 
wq[2][0] = -4; wq[2][1] = 8; wq[2][2] = -8; wq[2][3] = -15; wq[2][4] = -9; wq[2][5] = -16; wq[2][6] = 10; wq[2][7] = -13; wq[2][8] = 13; wq[2][9] = -14; wq[2][10] = 15; wq[2][11] = -8; wq[2][12] = -5; wq[2][13] = -16; wq[2][14] = -11; wq[2][15] = -10; 
wq[3][0] = 5; wq[3][1] = 11; wq[3][2] = -13; wq[3][3] = -3; wq[3][4] = -7; wq[3][5] = -7; wq[3][6] = -9; wq[3][7] = 13; wq[3][8] = -7; wq[3][9] = -7; wq[3][10] = 5; wq[3][11] = -7; wq[3][12] = 8; wq[3][13] = 1; wq[3][14] = 6; wq[3][15] = 4; 
wq[4][0] = -13; wq[4][1] = 5; wq[4][2] = -11; wq[4][3] = -14; wq[4][4] = 11; wq[4][5] = -11; wq[4][6] = 7; wq[4][7] = 3; wq[4][8] = 9; wq[4][9] = -7; wq[4][10] = 16; wq[4][11] = -4; wq[4][12] = -8; wq[4][13] = 13; wq[4][14] = -16; wq[4][15] = -6; 
wq[5][0] = -3; wq[5][1] = 3; wq[5][2] = -13; wq[5][3] = 6; wq[5][4] = 4; wq[5][5] = -13; wq[5][6] = 13; wq[5][7] = 10; wq[5][8] = -9; wq[5][9] = -12; wq[5][10] = -16; wq[5][11] = -11; wq[5][12] = 10; wq[5][13] = 9; wq[5][14] = 13; wq[5][15] = 3; 
wq[6][0] = -6; wq[6][1] = 15; wq[6][2] = 3; wq[6][3] = 16; wq[6][4] = 3; wq[6][5] = -2; wq[6][6] = -15; wq[6][7] = -6; wq[6][8] = -6; wq[6][9] = -6; wq[6][10] = -14; wq[6][11] = -14; wq[6][12] = 15; wq[6][13] = -15; wq[6][14] = 0; wq[6][15] = 0; 
wq[7][0] = -1; wq[7][1] = 14; wq[7][2] = 4; wq[7][3] = 2; wq[7][4] = -10; wq[7][5] = 15; wq[7][6] = 6; wq[7][7] = -4; wq[7][8] = -4; wq[7][9] = -14; wq[7][10] = 14; wq[7][11] = -9; wq[7][12] = -4; wq[7][13] = -13; wq[7][14] = -11; wq[7][15] = -5; 
wq[8][0] = 9; wq[8][1] = -2; wq[8][2] = -4; wq[8][3] = 14; wq[8][4] = -13; wq[8][5] = -11; wq[8][6] = 16; wq[8][7] = 4; wq[8][8] = 14; wq[8][9] = 9; wq[8][10] = -10; wq[8][11] = -1; wq[8][12] = -12; wq[8][13] = 1; wq[8][14] = 7; wq[8][15] = -8; 
wq[9][0] = 12; wq[9][1] = -15; wq[9][2] = 10; wq[9][3] = 13; wq[9][4] = -11; wq[9][5] = -7; wq[9][6] = -14; wq[9][7] = 12; wq[9][8] = 7; wq[9][9] = 13; wq[9][10] = -12; wq[9][11] = 6; wq[9][12] = 8; wq[9][13] = 11; wq[9][14] = 1; wq[9][15] = -6; 
wq[10][0] = 7; wq[10][1] = -6; wq[10][2] = -8; wq[10][3] = -6; wq[10][4] = 2; wq[10][5] = 7; wq[10][6] = -12; wq[10][7] = -12; wq[10][8] = 12; wq[10][9] = 2; wq[10][10] = 11; wq[10][11] = -13; wq[10][12] = 14; wq[10][13] = 15; wq[10][14] = 0; wq[10][15] = -2; 
wq[11][0] = 4; wq[11][1] = 5; wq[11][2] = -10; wq[11][3] = -1; wq[11][4] = -16; wq[11][5] = -6; wq[11][6] = -9; wq[11][7] = -16; wq[11][8] = -4; wq[11][9] = 14; wq[11][10] = 2; wq[11][11] = -10; wq[11][12] = 3; wq[11][13] = 8; wq[11][14] = 8; wq[11][15] = 11; 
wq[12][0] = -15; wq[12][1] = 9; wq[12][2] = 14; wq[12][3] = 5; wq[12][4] = -14; wq[12][5] = -16; wq[12][6] = 1; wq[12][7] = 15; wq[12][8] = 12; wq[12][9] = -3; wq[12][10] = 6; wq[12][11] = -7; wq[12][12] = -11; wq[12][13] = -12; wq[12][14] = 15; wq[12][15] = -13; 
wq[13][0] = -14; wq[13][1] = -11; wq[13][2] = -14; wq[13][3] = -8; wq[13][4] = 10; wq[13][5] = 3; wq[13][6] = 7; wq[13][7] = 2; wq[13][8] = 8; wq[13][9] = 13; wq[13][10] = 8; wq[13][11] = -14; wq[13][12] = 13; wq[13][13] = -6; wq[13][14] = 15; wq[13][15] = -2; 
wq[14][0] = 3; wq[14][1] = 2; wq[14][2] = -13; wq[14][3] = 1; wq[14][4] = -15; wq[14][5] = 9; wq[14][6] = -16; wq[14][7] = -4; wq[14][8] = 16; wq[14][9] = -10; wq[14][10] = -2; wq[14][11] = 3; wq[14][12] = -15; wq[14][13] = 8; wq[14][14] = -13; wq[14][15] = 7; 
wq[15][0] = -13; wq[15][1] = 10; wq[15][2] = 11; wq[15][3] = -9; wq[15][4] = -4; wq[15][5] = 0; wq[15][6] = -9; wq[15][7] = -1; wq[15][8] = 14; wq[15][9] = -4; wq[15][10] = 11; wq[15][11] = 0; wq[15][12] = -7; wq[15][13] = 9; wq[15][14] = 9; wq[15][15] = -13; 
wq[16][0] = -10; wq[16][1] = 1; wq[16][2] = -13; wq[16][3] = 9; wq[16][4] = -10; wq[16][5] = 3; wq[16][6] = 11; wq[16][7] = 12; wq[16][8] = -3; wq[16][9] = -12; wq[16][10] = 1; wq[16][11] = 6; wq[16][12] = -3; wq[16][13] = 15; wq[16][14] = 12; wq[16][15] = 4; 
wq[17][0] = 9; wq[17][1] = 15; wq[17][2] = -14; wq[17][3] = -14; wq[17][4] = -12; wq[17][5] = -6; wq[17][6] = -6; wq[17][7] = -1; wq[17][8] = -12; wq[17][9] = -10; wq[17][10] = -6; wq[17][11] = -12; wq[17][12] = -9; wq[17][13] = -13; wq[17][14] = 12; wq[17][15] = -10; 
wq[18][0] = 7; wq[18][1] = 4; wq[18][2] = -3; wq[18][3] = 12; wq[18][4] = 12; wq[18][5] = -16; wq[18][6] = -10; wq[18][7] = 3; wq[18][8] = 3; wq[18][9] = -7; wq[18][10] = 8; wq[18][11] = -1; wq[18][12] = 0; wq[18][13] = -12; wq[18][14] = 9; wq[18][15] = 2; 
wq[19][0] = -1; wq[19][1] = -5; wq[19][2] = -9; wq[19][3] = 14; wq[19][4] = -11; wq[19][5] = -10; wq[19][6] = 11; wq[19][7] = 6; wq[19][8] = 16; wq[19][9] = 16; wq[19][10] = -9; wq[19][11] = 8; wq[19][12] = -9; wq[19][13] = 6; wq[19][14] = -10; wq[19][15] = 5; 
wq[20][0] = -12; wq[20][1] = -9; wq[20][2] = 4; wq[20][3] = -14; wq[20][4] = 0; wq[20][5] = -7; wq[20][6] = 3; wq[20][7] = 13; wq[20][8] = -16; wq[20][9] = 16; wq[20][10] = -3; wq[20][11] = -12; wq[20][12] = 14; wq[20][13] = 12; wq[20][14] = 7; wq[20][15] = -14; 
wq[21][0] = 7; wq[21][1] = -8; wq[21][2] = 2; wq[21][3] = 11; wq[21][4] = 16; wq[21][5] = 12; wq[21][6] = -6; wq[21][7] = -14; wq[21][8] = -14; wq[21][9] = -3; wq[21][10] = 10; wq[21][11] = 10; wq[21][12] = 1; wq[21][13] = -2; wq[21][14] = -5; wq[21][15] = -4; 
wq[22][0] = 9; wq[22][1] = -12; wq[22][2] = -14; wq[22][3] = -13; wq[22][4] = 1; wq[22][5] = 5; wq[22][6] = 4; wq[22][7] = 12; wq[22][8] = 12; wq[22][9] = 1; wq[22][10] = -8; wq[22][11] = -1; wq[22][12] = -7; wq[22][13] = -10; wq[22][14] = -14; wq[22][15] = -10; 
wq[23][0] = -1; wq[23][1] = -12; wq[23][2] = -3; wq[23][3] = 16; wq[23][4] = 16; wq[23][5] = 15; wq[23][6] = 6; wq[23][7] = -8; wq[23][8] = -12; wq[23][9] = -12; wq[23][10] = 13; wq[23][11] = -12; wq[23][12] = -1; wq[23][13] = -6; wq[23][14] = 9; wq[23][15] = -7; 
wq[24][0] = 12; wq[24][1] = 9; wq[24][2] = -12; wq[24][3] = 9; wq[24][4] = -5; wq[24][5] = 8; wq[24][6] = 12; wq[24][7] = 12; wq[24][8] = -15; wq[24][9] = 14; wq[24][10] = -14; wq[24][11] = 12; wq[24][12] = 14; wq[24][13] = 3; wq[24][14] = 1; wq[24][15] = -6; 
wq[25][0] = 10; wq[25][1] = 3; wq[25][2] = 12; wq[25][3] = 6; wq[25][4] = 13; wq[25][5] = -4; wq[25][6] = -8; wq[25][7] = -4; wq[25][8] = 10; wq[25][9] = -14; wq[25][10] = 9; wq[25][11] = -5; wq[25][12] = 16; wq[25][13] = 16; wq[25][14] = 9; wq[25][15] = -13; 
wq[26][0] = 5; wq[26][1] = -12; wq[26][2] = 9; wq[26][3] = -8; wq[26][4] = -8; wq[26][5] = 15; wq[26][6] = -11; wq[26][7] = 7; wq[26][8] = -1; wq[26][9] = 7; wq[26][10] = -16; wq[26][11] = -1; wq[26][12] = -2; wq[26][13] = -4; wq[26][14] = -13; wq[26][15] = 0; 
wq[27][0] = 2; wq[27][1] = 14; wq[27][2] = 11; wq[27][3] = 1; wq[27][4] = 11; wq[27][5] = 12; wq[27][6] = 12; wq[27][7] = -9; wq[27][8] = 2; wq[27][9] = -4; wq[27][10] = -6; wq[27][11] = -16; wq[27][12] = 4; wq[27][13] = 8; wq[27][14] = 4; wq[27][15] = 2; 
wq[28][0] = 10; wq[28][1] = 6; wq[28][2] = -6; wq[28][3] = 9; wq[28][4] = 3; wq[28][5] = -11; wq[28][6] = 8; wq[28][7] = -9; wq[28][8] = 12; wq[28][9] = -6; wq[28][10] = 14; wq[28][11] = 12; wq[28][12] = -9; wq[28][13] = 12; wq[28][14] = 9; wq[28][15] = -5; 
wq[29][0] = 12; wq[29][1] = -5; wq[29][2] = -10; wq[29][3] = 2; wq[29][4] = 6; wq[29][5] = 14; wq[29][6] = 16; wq[29][7] = -7; wq[29][8] = -15; wq[29][9] = -5; wq[29][10] = 7; wq[29][11] = -13; wq[29][12] = 5; wq[29][13] = 5; wq[29][14] = 10; wq[29][15] = 0; 
wq[30][0] = 7; wq[30][1] = 1; wq[30][2] = -5; wq[30][3] = 15; wq[30][4] = -15; wq[30][5] = 9; wq[30][6] = 8; wq[30][7] = -13; wq[30][8] = 4; wq[30][9] = 7; wq[30][10] = -12; wq[30][11] = -4; wq[30][12] = -15; wq[30][13] = 5; wq[30][14] = 10; wq[30][15] = 13; 
wq[31][0] = -10; wq[31][1] = 9; wq[31][2] = -3; wq[31][3] = -5; wq[31][4] = 4; wq[31][5] = -15; wq[31][6] = 11; wq[31][7] = 0; wq[31][8] = -13; wq[31][9] = -14; wq[31][10] = 13; wq[31][11] = 2; wq[31][12] = -5; wq[31][13] = -16; wq[31][14] = -15; wq[31][15] = 16; 
wq[32][0] = 0; wq[32][1] = 7; wq[32][2] = 13; wq[32][3] = -10; wq[32][4] = 4; wq[32][5] = 16; wq[32][6] = 13; wq[32][7] = 13; wq[32][8] = -8; wq[32][9] = -14; wq[32][10] = 7; wq[32][11] = -4; wq[32][12] = -7; wq[32][13] = 10; wq[32][14] = -10; wq[32][15] = -15; 
wq[33][0] = 11; wq[33][1] = -2; wq[33][2] = 1; wq[33][3] = 7; wq[33][4] = -11; wq[33][5] = 15; wq[33][6] = -3; wq[33][7] = -11; wq[33][8] = 9; wq[33][9] = -4; wq[33][10] = -2; wq[33][11] = 16; wq[33][12] = -5; wq[33][13] = -4; wq[33][14] = -9; wq[33][15] = 6; 
wq[34][0] = -6; wq[34][1] = -8; wq[34][2] = 0; wq[34][3] = 10; wq[34][4] = -8; wq[34][5] = 7; wq[34][6] = -2; wq[34][7] = -2; wq[34][8] = 2; wq[34][9] = -9; wq[34][10] = 12; wq[34][11] = -13; wq[34][12] = -13; wq[34][13] = -4; wq[34][14] = -16; wq[34][15] = 15; 
wq[35][0] = 1; wq[35][1] = -13; wq[35][2] = -10; wq[35][3] = 8; wq[35][4] = -12; wq[35][5] = -9; wq[35][6] = -13; wq[35][7] = 11; wq[35][8] = -8; wq[35][9] = -10; wq[35][10] = 7; wq[35][11] = 10; wq[35][12] = 0; wq[35][13] = -16; wq[35][14] = 13; wq[35][15] = 8; 
wq[36][0] = 7; wq[36][1] = -16; wq[36][2] = 3; wq[36][3] = -10; wq[36][4] = 15; wq[36][5] = -4; wq[36][6] = 13; wq[36][7] = 9; wq[36][8] = 0; wq[36][9] = 2; wq[36][10] = -9; wq[36][11] = -3; wq[36][12] = -6; wq[36][13] = 12; wq[36][14] = 3; wq[36][15] = 12; 
wq[37][0] = -8; wq[37][1] = 16; wq[37][2] = 11; wq[37][3] = 1; wq[37][4] = -16; wq[37][5] = -14; wq[37][6] = -12; wq[37][7] = -4; wq[37][8] = -1; wq[37][9] = 12; wq[37][10] = -13; wq[37][11] = -8; wq[37][12] = 1; wq[37][13] = 12; wq[37][14] = 7; wq[37][15] = 3; 
wq[38][0] = 16; wq[38][1] = 1; wq[38][2] = 7; wq[38][3] = -12; wq[38][4] = 0; wq[38][5] = 0; wq[38][6] = -10; wq[38][7] = 10; wq[38][8] = -5; wq[38][9] = -1; wq[38][10] = 16; wq[38][11] = -6; wq[38][12] = 1; wq[38][13] = -16; wq[38][14] = -10; wq[38][15] = 10; 
wq[39][0] = 0; wq[39][1] = 5; wq[39][2] = 13; wq[39][3] = 14; wq[39][4] = 7; wq[39][5] = 16; wq[39][6] = -16; wq[39][7] = -2; wq[39][8] = -15; wq[39][9] = -14; wq[39][10] = -2; wq[39][11] = -6; wq[39][12] = -13; wq[39][13] = 10; wq[39][14] = 4; wq[39][15] = 7; 
wq[40][0] = 2; wq[40][1] = 15; wq[40][2] = -9; wq[40][3] = -2; wq[40][4] = 9; wq[40][5] = -10; wq[40][6] = -11; wq[40][7] = 14; wq[40][8] = 14; wq[40][9] = 10; wq[40][10] = 1; wq[40][11] = 16; wq[40][12] = 15; wq[40][13] = -2; wq[40][14] = -5; wq[40][15] = 9; 
wq[41][0] = -12; wq[41][1] = -11; wq[41][2] = 5; wq[41][3] = 16; wq[41][4] = 15; wq[41][5] = 8; wq[41][6] = -8; wq[41][7] = 7; wq[41][8] = -6; wq[41][9] = 9; wq[41][10] = -15; wq[41][11] = 13; wq[41][12] = 10; wq[41][13] = 9; wq[41][14] = -1; wq[41][15] = 10; 
wq[42][0] = -9; wq[42][1] = 16; wq[42][2] = 7; wq[42][3] = 4; wq[42][4] = -9; wq[42][5] = 1; wq[42][6] = -3; wq[42][7] = -13; wq[42][8] = -7; wq[42][9] = 16; wq[42][10] = 10; wq[42][11] = -3; wq[42][12] = -9; wq[42][13] = 12; wq[42][14] = 14; wq[42][15] = -8; 
wq[43][0] = -6; wq[43][1] = 6; wq[43][2] = 2; wq[43][3] = -8; wq[43][4] = -10; wq[43][5] = -2; wq[43][6] = -5; wq[43][7] = -8; wq[43][8] = -8; wq[43][9] = -12; wq[43][10] = 13; wq[43][11] = 7; wq[43][12] = 4; wq[43][13] = 0; wq[43][14] = 10; wq[43][15] = -4; 
wq[44][0] = 2; wq[44][1] = -10; wq[44][2] = 4; wq[44][3] = -16; wq[44][4] = 11; wq[44][5] = 7; wq[44][6] = -4; wq[44][7] = -11; wq[44][8] = -14; wq[44][9] = 15; wq[44][10] = 2; wq[44][11] = -7; wq[44][12] = 2; wq[44][13] = 10; wq[44][14] = -15; wq[44][15] = 15; 
wq[45][0] = 12; wq[45][1] = 15; wq[45][2] = 10; wq[45][3] = -5; wq[45][4] = 0; wq[45][5] = -10; wq[45][6] = -15; wq[45][7] = -13; wq[45][8] = -14; wq[45][9] = 1; wq[45][10] = -3; wq[45][11] = -7; wq[45][12] = -6; wq[45][13] = 7; wq[45][14] = -14; wq[45][15] = 15; 
wq[46][0] = -10; wq[46][1] = -13; wq[46][2] = 13; wq[46][3] = 11; wq[46][4] = -11; wq[46][5] = 3; wq[46][6] = 14; wq[46][7] = 1; wq[46][8] = 14; wq[46][9] = -2; wq[46][10] = 3; wq[46][11] = 11; wq[46][12] = 13; wq[46][13] = 15; wq[46][14] = 5; wq[46][15] = 11; 
wq[47][0] = 3; wq[47][1] = -3; wq[47][2] = 4; wq[47][3] = -3; wq[47][4] = 11; wq[47][5] = -1; wq[47][6] = -6; wq[47][7] = -8; wq[47][8] = 13; wq[47][9] = -3; wq[47][10] = 13; wq[47][11] = 0; wq[47][12] = -10; wq[47][13] = 12; wq[47][14] = -12; wq[47][15] = 9; 
wq[48][0] = 5; wq[48][1] = 5; wq[48][2] = -7; wq[48][3] = -3; wq[48][4] = -2; wq[48][5] = -11; wq[48][6] = -14; wq[48][7] = 2; wq[48][8] = 13; wq[48][9] = 10; wq[48][10] = -4; wq[48][11] = -2; wq[48][12] = 9; wq[48][13] = 14; wq[48][14] = -11; wq[48][15] = -11; 
wq[49][0] = 15; wq[49][1] = -10; wq[49][2] = -11; wq[49][3] = 7; wq[49][4] = -13; wq[49][5] = -15; wq[49][6] = -9; wq[49][7] = 10; wq[49][8] = 14; wq[49][9] = -10; wq[49][10] = 6; wq[49][11] = 9; wq[49][12] = 14; wq[49][13] = 8; wq[49][14] = 0; wq[49][15] = -11; 
wq[50][0] = 4; wq[50][1] = 10; wq[50][2] = 7; wq[50][3] = -13; wq[50][4] = 9; wq[50][5] = -7; wq[50][6] = -11; wq[50][7] = -16; wq[50][8] = 1; wq[50][9] = -7; wq[50][10] = 8; wq[50][11] = -12; wq[50][12] = 11; wq[50][13] = 10; wq[50][14] = 4; wq[50][15] = -1; 
wq[51][0] = -8; wq[51][1] = 11; wq[51][2] = -14; wq[51][3] = -5; wq[51][4] = -11; wq[51][5] = -10; wq[51][6] = 3; wq[51][7] = -8; wq[51][8] = 4; wq[51][9] = -3; wq[51][10] = -15; wq[51][11] = 8; wq[51][12] = -6; wq[51][13] = -5; wq[51][14] = 5; wq[51][15] = 2; 
wq[52][0] = 16; wq[52][1] = 4; wq[52][2] = -7; wq[52][3] = 6; wq[52][4] = -8; wq[52][5] = -7; wq[52][6] = 2; wq[52][7] = 12; wq[52][8] = 1; wq[52][9] = -4; wq[52][10] = -6; wq[52][11] = 3; wq[52][12] = -9; wq[52][13] = 16; wq[52][14] = -5; wq[52][15] = -7; 
wq[53][0] = -11; wq[53][1] = -6; wq[53][2] = -16; wq[53][3] = 14; wq[53][4] = 5; wq[53][5] = 0; wq[53][6] = -8; wq[53][7] = -4; wq[53][8] = 4; wq[53][9] = 3; wq[53][10] = -16; wq[53][11] = -1; wq[53][12] = -2; wq[53][13] = -4; wq[53][14] = 14; wq[53][15] = -12; 
wq[54][0] = -1; wq[54][1] = 0; wq[54][2] = 6; wq[54][3] = -4; wq[54][4] = 3; wq[54][5] = -4; wq[54][6] = 9; wq[54][7] = 10; wq[54][8] = 1; wq[54][9] = 0; wq[54][10] = -6; wq[54][11] = 14; wq[54][12] = 10; wq[54][13] = -16; wq[54][14] = 0; wq[54][15] = -12; 
wq[55][0] = -14; wq[55][1] = -7; wq[55][2] = 6; wq[55][3] = -7; wq[55][4] = -2; wq[55][5] = 4; wq[55][6] = 16; wq[55][7] = 14; wq[55][8] = 14; wq[55][9] = 2; wq[55][10] = 1; wq[55][11] = 2; wq[55][12] = -16; wq[55][13] = 1; wq[55][14] = -5; wq[55][15] = -11; 
wq[56][0] = -6; wq[56][1] = 10; wq[56][2] = 6; wq[56][3] = -1; wq[56][4] = 10; wq[56][5] = 7; wq[56][6] = -4; wq[56][7] = 10; wq[56][8] = 3; wq[56][9] = -3; wq[56][10] = -4; wq[56][11] = 13; wq[56][12] = -10; wq[56][13] = -5; wq[56][14] = 10; wq[56][15] = 9; 
wq[57][0] = -15; wq[57][1] = 2; wq[57][2] = 14; wq[57][3] = -8; wq[57][4] = -6; wq[57][5] = -10; wq[57][6] = 6; wq[57][7] = -14; wq[57][8] = 7; wq[57][9] = 14; wq[57][10] = -14; wq[57][11] = 3; wq[57][12] = -12; wq[57][13] = 8; wq[57][14] = 10; wq[57][15] = -4; 
wq[58][0] = -16; wq[58][1] = 8; wq[58][2] = 7; wq[58][3] = 7; wq[58][4] = -3; wq[58][5] = -4; wq[58][6] = -10; wq[58][7] = 4; wq[58][8] = 15; wq[58][9] = 15; wq[58][10] = -8; wq[58][11] = 9; wq[58][12] = -4; wq[58][13] = -9; wq[58][14] = 8; wq[58][15] = -2; 
wq[59][0] = -14; wq[59][1] = -3; wq[59][2] = -13; wq[59][3] = 5; wq[59][4] = 12; wq[59][5] = 12; wq[59][6] = 7; wq[59][7] = 11; wq[59][8] = 7; wq[59][9] = -2; wq[59][10] = 10; wq[59][11] = -13; wq[59][12] = -16; wq[59][13] = -15; wq[59][14] = -3; wq[59][15] = 16; 
wq[60][0] = 12; wq[60][1] = 2; wq[60][2] = -4; wq[60][3] = -12; wq[60][4] = -10; wq[60][5] = 16; wq[60][6] = 5; wq[60][7] = -3; wq[60][8] = 14; wq[60][9] = 14; wq[60][10] = 11; wq[60][11] = 7; wq[60][12] = 4; wq[60][13] = 0; wq[60][14] = 11; wq[60][15] = 3; 
wq[61][0] = 6; wq[61][1] = 15; wq[61][2] = -10; wq[61][3] = -5; wq[61][4] = -16; wq[61][5] = 3; wq[61][6] = -10; wq[61][7] = -12; wq[61][8] = 14; wq[61][9] = 1; wq[61][10] = 1; wq[61][11] = -4; wq[61][12] = -10; wq[61][13] = 3; wq[61][14] = -2; wq[61][15] = -14; 
wq[62][0] = 7; wq[62][1] = 16; wq[62][2] = 13; wq[62][3] = 0; wq[62][4] = 4; wq[62][5] = -4; wq[62][6] = 8; wq[62][7] = -6; wq[62][8] = 6; wq[62][9] = 1; wq[62][10] = -3; wq[62][11] = -9; wq[62][12] = 15; wq[62][13] = 1; wq[62][14] = 15; wq[62][15] = 8; 
wq[63][0] = 16; wq[63][1] = 4; wq[63][2] = -13; wq[63][3] = 11; wq[63][4] = -14; wq[63][5] = -12; wq[63][6] = 5; wq[63][7] = -7; wq[63][8] = 9; wq[63][9] = 16; wq[63][10] = -3; wq[63][11] = 11; wq[63][12] = -16; wq[63][13] = -11; wq[63][14] = 7; wq[63][15] = -12; 

wk[0][0] = 12; wk[0][1] = 12; wk[0][2] = 11; wk[0][3] = 13; wk[0][4] = -10; wk[0][5] = -14; wk[0][6] = 11; wk[0][7] = -13; wk[0][8] = 3; wk[0][9] = -5; wk[0][10] = -5; wk[0][11] = 9; wk[0][12] = 6; wk[0][13] = -6; wk[0][14] = 13; wk[0][15] = -5; 
wk[1][0] = -7; wk[1][1] = -10; wk[1][2] = -1; wk[1][3] = 3; wk[1][4] = 6; wk[1][5] = 2; wk[1][6] = 8; wk[1][7] = 16; wk[1][8] = 9; wk[1][9] = 6; wk[1][10] = -15; wk[1][11] = -14; wk[1][12] = 5; wk[1][13] = 6; wk[1][14] = -6; wk[1][15] = -8; 
wk[2][0] = -1; wk[2][1] = 10; wk[2][2] = -16; wk[2][3] = -13; wk[2][4] = 8; wk[2][5] = 11; wk[2][6] = -13; wk[2][7] = 8; wk[2][8] = 5; wk[2][9] = 9; wk[2][10] = 7; wk[2][11] = 0; wk[2][12] = -11; wk[2][13] = -7; wk[2][14] = 3; wk[2][15] = -9; 
wk[3][0] = -16; wk[3][1] = 16; wk[3][2] = -13; wk[3][3] = -16; wk[3][4] = 3; wk[3][5] = -15; wk[3][6] = 14; wk[3][7] = 13; wk[3][8] = -15; wk[3][9] = 12; wk[3][10] = 16; wk[3][11] = -14; wk[3][12] = -6; wk[3][13] = -3; wk[3][14] = 8; wk[3][15] = 4; 
wk[4][0] = 13; wk[4][1] = -13; wk[4][2] = -14; wk[4][3] = -16; wk[4][4] = -2; wk[4][5] = -10; wk[4][6] = 13; wk[4][7] = -5; wk[4][8] = -4; wk[4][9] = 8; wk[4][10] = 15; wk[4][11] = -12; wk[4][12] = -12; wk[4][13] = -11; wk[4][14] = 13; wk[4][15] = 7; 
wk[5][0] = -1; wk[5][1] = 0; wk[5][2] = 15; wk[5][3] = 5; wk[5][4] = 2; wk[5][5] = 10; wk[5][6] = -6; wk[5][7] = 11; wk[5][8] = 13; wk[5][9] = 8; wk[5][10] = 0; wk[5][11] = 10; wk[5][12] = 14; wk[5][13] = -15; wk[5][14] = 15; wk[5][15] = -7; 
wk[6][0] = -2; wk[6][1] = 13; wk[6][2] = 12; wk[6][3] = 7; wk[6][4] = -5; wk[6][5] = 7; wk[6][6] = -14; wk[6][7] = 10; wk[6][8] = -4; wk[6][9] = 13; wk[6][10] = 16; wk[6][11] = -15; wk[6][12] = 13; wk[6][13] = 10; wk[6][14] = -15; wk[6][15] = -14; 
wk[7][0] = -9; wk[7][1] = 2; wk[7][2] = 11; wk[7][3] = 11; wk[7][4] = 14; wk[7][5] = 11; wk[7][6] = -12; wk[7][7] = 4; wk[7][8] = -16; wk[7][9] = -6; wk[7][10] = 7; wk[7][11] = 8; wk[7][12] = -12; wk[7][13] = 0; wk[7][14] = -11; wk[7][15] = -6; 
wk[8][0] = -4; wk[8][1] = 11; wk[8][2] = -2; wk[8][3] = -8; wk[8][4] = -5; wk[8][5] = 9; wk[8][6] = -2; wk[8][7] = 15; wk[8][8] = -1; wk[8][9] = 13; wk[8][10] = 10; wk[8][11] = -13; wk[8][12] = 1; wk[8][13] = 5; wk[8][14] = -8; wk[8][15] = -12; 
wk[9][0] = -9; wk[9][1] = -6; wk[9][2] = -1; wk[9][3] = -12; wk[9][4] = 5; wk[9][5] = -13; wk[9][6] = -13; wk[9][7] = 10; wk[9][8] = 2; wk[9][9] = 5; wk[9][10] = 0; wk[9][11] = -10; wk[9][12] = 4; wk[9][13] = 9; wk[9][14] = -9; wk[9][15] = -16; 
wk[10][0] = 11; wk[10][1] = 4; wk[10][2] = -13; wk[10][3] = -7; wk[10][4] = 6; wk[10][5] = 3; wk[10][6] = -4; wk[10][7] = -12; wk[10][8] = -1; wk[10][9] = -13; wk[10][10] = 5; wk[10][11] = 7; wk[10][12] = 15; wk[10][13] = -16; wk[10][14] = 14; wk[10][15] = 8; 
wk[11][0] = 1; wk[11][1] = -9; wk[11][2] = 0; wk[11][3] = -5; wk[11][4] = 16; wk[11][5] = 5; wk[11][6] = -6; wk[11][7] = 5; wk[11][8] = 12; wk[11][9] = -8; wk[11][10] = 16; wk[11][11] = -7; wk[11][12] = 3; wk[11][13] = -6; wk[11][14] = -16; wk[11][15] = 10; 
wk[12][0] = -6; wk[12][1] = -4; wk[12][2] = 8; wk[12][3] = -2; wk[12][4] = -16; wk[12][5] = -8; wk[12][6] = -1; wk[12][7] = 10; wk[12][8] = 7; wk[12][9] = -5; wk[12][10] = -15; wk[12][11] = 15; wk[12][12] = -8; wk[12][13] = 3; wk[12][14] = 14; wk[12][15] = 14; 
wk[13][0] = 7; wk[13][1] = 6; wk[13][2] = -9; wk[13][3] = -14; wk[13][4] = -13; wk[13][5] = -14; wk[13][6] = 5; wk[13][7] = 8; wk[13][8] = -16; wk[13][9] = -2; wk[13][10] = 6; wk[13][11] = -13; wk[13][12] = 3; wk[13][13] = -6; wk[13][14] = -10; wk[13][15] = 4; 
wk[14][0] = -16; wk[14][1] = -9; wk[14][2] = -8; wk[14][3] = -2; wk[14][4] = 3; wk[14][5] = 12; wk[14][6] = -8; wk[14][7] = 6; wk[14][8] = 2; wk[14][9] = 12; wk[14][10] = 8; wk[14][11] = -1; wk[14][12] = -12; wk[14][13] = -3; wk[14][14] = -11; wk[14][15] = -10; 
wk[15][0] = -12; wk[15][1] = -1; wk[15][2] = 15; wk[15][3] = -15; wk[15][4] = -12; wk[15][5] = -12; wk[15][6] = 3; wk[15][7] = 12; wk[15][8] = 4; wk[15][9] = 11; wk[15][10] = -8; wk[15][11] = -7; wk[15][12] = 2; wk[15][13] = -3; wk[15][14] = -10; wk[15][15] = -6; 
wk[16][0] = -7; wk[16][1] = -2; wk[16][2] = -13; wk[16][3] = 16; wk[16][4] = -8; wk[16][5] = -13; wk[16][6] = 4; wk[16][7] = 11; wk[16][8] = -6; wk[16][9] = -14; wk[16][10] = 4; wk[16][11] = -13; wk[16][12] = 9; wk[16][13] = 11; wk[16][14] = 6; wk[16][15] = -2; 
wk[17][0] = -14; wk[17][1] = 13; wk[17][2] = 12; wk[17][3] = 14; wk[17][4] = -1; wk[17][5] = -3; wk[17][6] = -13; wk[17][7] = -7; wk[17][8] = -1; wk[17][9] = -13; wk[17][10] = -8; wk[17][11] = 13; wk[17][12] = -10; wk[17][13] = -10; wk[17][14] = -12; wk[17][15] = -4; 
wk[18][0] = -6; wk[18][1] = -4; wk[18][2] = 11; wk[18][3] = 13; wk[18][4] = -16; wk[18][5] = 0; wk[18][6] = 10; wk[18][7] = 11; wk[18][8] = -6; wk[18][9] = -9; wk[18][10] = 1; wk[18][11] = -14; wk[18][12] = 11; wk[18][13] = 0; wk[18][14] = -1; wk[18][15] = -2; 
wk[19][0] = -15; wk[19][1] = -4; wk[19][2] = 0; wk[19][3] = -9; wk[19][4] = 9; wk[19][5] = 9; wk[19][6] = 10; wk[19][7] = 5; wk[19][8] = -10; wk[19][9] = -13; wk[19][10] = 15; wk[19][11] = -12; wk[19][12] = -8; wk[19][13] = 3; wk[19][14] = 11; wk[19][15] = -3; 
wk[20][0] = 11; wk[20][1] = 13; wk[20][2] = 5; wk[20][3] = -15; wk[20][4] = 11; wk[20][5] = -8; wk[20][6] = -13; wk[20][7] = 7; wk[20][8] = 2; wk[20][9] = 1; wk[20][10] = 16; wk[20][11] = -4; wk[20][12] = 5; wk[20][13] = 5; wk[20][14] = -6; wk[20][15] = 0; 
wk[21][0] = 3; wk[21][1] = 13; wk[21][2] = 0; wk[21][3] = -12; wk[21][4] = 6; wk[21][5] = 6; wk[21][6] = 7; wk[21][7] = -3; wk[21][8] = -10; wk[21][9] = 5; wk[21][10] = -16; wk[21][11] = -16; wk[21][12] = 8; wk[21][13] = 11; wk[21][14] = -14; wk[21][15] = 5; 
wk[22][0] = 14; wk[22][1] = -11; wk[22][2] = -2; wk[22][3] = 10; wk[22][4] = 13; wk[22][5] = -12; wk[22][6] = 14; wk[22][7] = 11; wk[22][8] = -1; wk[22][9] = -7; wk[22][10] = -15; wk[22][11] = -14; wk[22][12] = -11; wk[22][13] = 12; wk[22][14] = 15; wk[22][15] = -13; 
wk[23][0] = 8; wk[23][1] = 10; wk[23][2] = 14; wk[23][3] = 6; wk[23][4] = 11; wk[23][5] = 5; wk[23][6] = -12; wk[23][7] = 2; wk[23][8] = 3; wk[23][9] = 11; wk[23][10] = 8; wk[23][11] = 10; wk[23][12] = -6; wk[23][13] = -1; wk[23][14] = 9; wk[23][15] = 12; 
wk[24][0] = 10; wk[24][1] = -14; wk[24][2] = -11; wk[24][3] = 11; wk[24][4] = 9; wk[24][5] = 16; wk[24][6] = -7; wk[24][7] = -9; wk[24][8] = 9; wk[24][9] = 13; wk[24][10] = -1; wk[24][11] = -8; wk[24][12] = 12; wk[24][13] = 3; wk[24][14] = 15; wk[24][15] = 1; 
wk[25][0] = 4; wk[25][1] = 10; wk[25][2] = -9; wk[25][3] = -2; wk[25][4] = -10; wk[25][5] = 16; wk[25][6] = 1; wk[25][7] = 6; wk[25][8] = -3; wk[25][9] = 11; wk[25][10] = -15; wk[25][11] = 5; wk[25][12] = -14; wk[25][13] = -16; wk[25][14] = -15; wk[25][15] = -11; 
wk[26][0] = 1; wk[26][1] = 1; wk[26][2] = -9; wk[26][3] = -6; wk[26][4] = 8; wk[26][5] = 4; wk[26][6] = 8; wk[26][7] = 4; wk[26][8] = -9; wk[26][9] = 16; wk[26][10] = 15; wk[26][11] = 11; wk[26][12] = 8; wk[26][13] = 8; wk[26][14] = 14; wk[26][15] = 1; 
wk[27][0] = 8; wk[27][1] = 14; wk[27][2] = -15; wk[27][3] = -5; wk[27][4] = -9; wk[27][5] = 5; wk[27][6] = -13; wk[27][7] = 9; wk[27][8] = -2; wk[27][9] = 6; wk[27][10] = -16; wk[27][11] = -4; wk[27][12] = 5; wk[27][13] = -10; wk[27][14] = 1; wk[27][15] = 4; 
wk[28][0] = -14; wk[28][1] = 13; wk[28][2] = 3; wk[28][3] = -16; wk[28][4] = -15; wk[28][5] = 8; wk[28][6] = 1; wk[28][7] = -14; wk[28][8] = 15; wk[28][9] = -6; wk[28][10] = -7; wk[28][11] = -2; wk[28][12] = -11; wk[28][13] = -4; wk[28][14] = 14; wk[28][15] = -6; 
wk[29][0] = 0; wk[29][1] = 7; wk[29][2] = -7; wk[29][3] = 3; wk[29][4] = -4; wk[29][5] = -13; wk[29][6] = -14; wk[29][7] = 6; wk[29][8] = 9; wk[29][9] = 9; wk[29][10] = -8; wk[29][11] = -11; wk[29][12] = -6; wk[29][13] = -14; wk[29][14] = 7; wk[29][15] = -5; 
wk[30][0] = 4; wk[30][1] = 14; wk[30][2] = 6; wk[30][3] = 11; wk[30][4] = 8; wk[30][5] = 5; wk[30][6] = 5; wk[30][7] = -4; wk[30][8] = 4; wk[30][9] = 12; wk[30][10] = -9; wk[30][11] = 16; wk[30][12] = -5; wk[30][13] = 11; wk[30][14] = 0; wk[30][15] = -6; 
wk[31][0] = 6; wk[31][1] = 0; wk[31][2] = -16; wk[31][3] = -1; wk[31][4] = 12; wk[31][5] = 15; wk[31][6] = 6; wk[31][7] = -3; wk[31][8] = -12; wk[31][9] = -8; wk[31][10] = -9; wk[31][11] = 13; wk[31][12] = -14; wk[31][13] = -2; wk[31][14] = 9; wk[31][15] = -16; 
wk[32][0] = -1; wk[32][1] = -6; wk[32][2] = 10; wk[32][3] = -13; wk[32][4] = -13; wk[32][5] = 5; wk[32][6] = -2; wk[32][7] = 13; wk[32][8] = 0; wk[32][9] = -15; wk[32][10] = 12; wk[32][11] = -12; wk[32][12] = -7; wk[32][13] = -12; wk[32][14] = 13; wk[32][15] = -6; 
wk[33][0] = -5; wk[33][1] = 0; wk[33][2] = -4; wk[33][3] = -2; wk[33][4] = -8; wk[33][5] = -15; wk[33][6] = 10; wk[33][7] = 10; wk[33][8] = -11; wk[33][9] = 8; wk[33][10] = -13; wk[33][11] = 13; wk[33][12] = -10; wk[33][13] = -5; wk[33][14] = -5; wk[33][15] = 16; 
wk[34][0] = -13; wk[34][1] = -8; wk[34][2] = -2; wk[34][3] = 14; wk[34][4] = 15; wk[34][5] = -13; wk[34][6] = -9; wk[34][7] = 8; wk[34][8] = 11; wk[34][9] = 4; wk[34][10] = -11; wk[34][11] = 1; wk[34][12] = 12; wk[34][13] = -4; wk[34][14] = -12; wk[34][15] = 16; 
wk[35][0] = -12; wk[35][1] = -8; wk[35][2] = 8; wk[35][3] = 4; wk[35][4] = -11; wk[35][5] = 9; wk[35][6] = 6; wk[35][7] = 12; wk[35][8] = -3; wk[35][9] = 12; wk[35][10] = -12; wk[35][11] = 14; wk[35][12] = -3; wk[35][13] = 3; wk[35][14] = -9; wk[35][15] = -13; 
wk[36][0] = 9; wk[36][1] = -8; wk[36][2] = -6; wk[36][3] = 6; wk[36][4] = 4; wk[36][5] = -10; wk[36][6] = 12; wk[36][7] = 1; wk[36][8] = 8; wk[36][9] = 4; wk[36][10] = -1; wk[36][11] = -5; wk[36][12] = -6; wk[36][13] = 4; wk[36][14] = 15; wk[36][15] = -8; 
wk[37][0] = -15; wk[37][1] = 15; wk[37][2] = 2; wk[37][3] = 16; wk[37][4] = -6; wk[37][5] = 9; wk[37][6] = -10; wk[37][7] = -4; wk[37][8] = 9; wk[37][9] = 5; wk[37][10] = 11; wk[37][11] = 6; wk[37][12] = -5; wk[37][13] = 6; wk[37][14] = -7; wk[37][15] = -8; 
wk[38][0] = 11; wk[38][1] = 15; wk[38][2] = -2; wk[38][3] = -15; wk[38][4] = -12; wk[38][5] = -10; wk[38][6] = -4; wk[38][7] = -12; wk[38][8] = 4; wk[38][9] = 5; wk[38][10] = 5; wk[38][11] = 1; wk[38][12] = -11; wk[38][13] = 16; wk[38][14] = -12; wk[38][15] = -1; 
wk[39][0] = -6; wk[39][1] = 11; wk[39][2] = -12; wk[39][3] = 9; wk[39][4] = -2; wk[39][5] = -8; wk[39][6] = -7; wk[39][7] = 0; wk[39][8] = 4; wk[39][9] = -16; wk[39][10] = 5; wk[39][11] = -4; wk[39][12] = -8; wk[39][13] = 6; wk[39][14] = 13; wk[39][15] = -9; 
wk[40][0] = 9; wk[40][1] = -6; wk[40][2] = 1; wk[40][3] = -8; wk[40][4] = -1; wk[40][5] = -5; wk[40][6] = -1; wk[40][7] = -13; wk[40][8] = -14; wk[40][9] = -4; wk[40][10] = -4; wk[40][11] = 14; wk[40][12] = -2; wk[40][13] = -11; wk[40][14] = 14; wk[40][15] = -14; 
wk[41][0] = 9; wk[41][1] = 0; wk[41][2] = -4; wk[41][3] = -5; wk[41][4] = 14; wk[41][5] = 5; wk[41][6] = 0; wk[41][7] = 1; wk[41][8] = -11; wk[41][9] = 9; wk[41][10] = 10; wk[41][11] = -16; wk[41][12] = 9; wk[41][13] = -14; wk[41][14] = -14; wk[41][15] = 16; 
wk[42][0] = 14; wk[42][1] = -3; wk[42][2] = 4; wk[42][3] = 16; wk[42][4] = 12; wk[42][5] = 0; wk[42][6] = 11; wk[42][7] = -11; wk[42][8] = 7; wk[42][9] = 6; wk[42][10] = -3; wk[42][11] = 3; wk[42][12] = 15; wk[42][13] = -14; wk[42][14] = 10; wk[42][15] = -14; 
wk[43][0] = -8; wk[43][1] = -9; wk[43][2] = 0; wk[43][3] = 13; wk[43][4] = 11; wk[43][5] = 11; wk[43][6] = 6; wk[43][7] = 11; wk[43][8] = 10; wk[43][9] = -15; wk[43][10] = 14; wk[43][11] = 7; wk[43][12] = 5; wk[43][13] = 4; wk[43][14] = -4; wk[43][15] = -14; 
wk[44][0] = -2; wk[44][1] = -12; wk[44][2] = 5; wk[44][3] = -8; wk[44][4] = -7; wk[44][5] = -12; wk[44][6] = -9; wk[44][7] = -14; wk[44][8] = 13; wk[44][9] = 13; wk[44][10] = 15; wk[44][11] = -11; wk[44][12] = -15; wk[44][13] = -10; wk[44][14] = -3; wk[44][15] = -7; 
wk[45][0] = 3; wk[45][1] = 1; wk[45][2] = 1; wk[45][3] = -11; wk[45][4] = 3; wk[45][5] = 12; wk[45][6] = -2; wk[45][7] = -3; wk[45][8] = -9; wk[45][9] = -6; wk[45][10] = 3; wk[45][11] = 16; wk[45][12] = -8; wk[45][13] = -7; wk[45][14] = 0; wk[45][15] = -5; 
wk[46][0] = -8; wk[46][1] = -12; wk[46][2] = -3; wk[46][3] = -10; wk[46][4] = -11; wk[46][5] = 0; wk[46][6] = 10; wk[46][7] = 10; wk[46][8] = -8; wk[46][9] = 8; wk[46][10] = 10; wk[46][11] = 7; wk[46][12] = 15; wk[46][13] = 9; wk[46][14] = -2; wk[46][15] = 0; 
wk[47][0] = -6; wk[47][1] = 11; wk[47][2] = -9; wk[47][3] = 15; wk[47][4] = -15; wk[47][5] = -3; wk[47][6] = -6; wk[47][7] = -15; wk[47][8] = -9; wk[47][9] = 2; wk[47][10] = 16; wk[47][11] = 2; wk[47][12] = -1; wk[47][13] = 8; wk[47][14] = 10; wk[47][15] = 6; 
wk[48][0] = -5; wk[48][1] = 4; wk[48][2] = 10; wk[48][3] = 2; wk[48][4] = 4; wk[48][5] = -3; wk[48][6] = 9; wk[48][7] = 14; wk[48][8] = 8; wk[48][9] = 11; wk[48][10] = -1; wk[48][11] = 10; wk[48][12] = 10; wk[48][13] = -5; wk[48][14] = 7; wk[48][15] = -16; 
wk[49][0] = -12; wk[49][1] = -13; wk[49][2] = 13; wk[49][3] = 9; wk[49][4] = 13; wk[49][5] = -4; wk[49][6] = -3; wk[49][7] = 10; wk[49][8] = 8; wk[49][9] = -9; wk[49][10] = -7; wk[49][11] = 16; wk[49][12] = 3; wk[49][13] = 3; wk[49][14] = -3; wk[49][15] = -8; 
wk[50][0] = 10; wk[50][1] = 2; wk[50][2] = 8; wk[50][3] = 3; wk[50][4] = -4; wk[50][5] = -11; wk[50][6] = 13; wk[50][7] = -6; wk[50][8] = 1; wk[50][9] = 7; wk[50][10] = 12; wk[50][11] = 8; wk[50][12] = -11; wk[50][13] = -15; wk[50][14] = 11; wk[50][15] = 1; 
wk[51][0] = -14; wk[51][1] = 10; wk[51][2] = -16; wk[51][3] = 7; wk[51][4] = 16; wk[51][5] = -8; wk[51][6] = 4; wk[51][7] = -3; wk[51][8] = -9; wk[51][9] = 4; wk[51][10] = 15; wk[51][11] = -3; wk[51][12] = -6; wk[51][13] = -2; wk[51][14] = 5; wk[51][15] = 9; 
wk[52][0] = 1; wk[52][1] = -13; wk[52][2] = -4; wk[52][3] = -8; wk[52][4] = -4; wk[52][5] = 10; wk[52][6] = -11; wk[52][7] = -6; wk[52][8] = -2; wk[52][9] = -9; wk[52][10] = 2; wk[52][11] = 9; wk[52][12] = -15; wk[52][13] = 12; wk[52][14] = -15; wk[52][15] = 10; 
wk[53][0] = 12; wk[53][1] = 1; wk[53][2] = 13; wk[53][3] = 0; wk[53][4] = 1; wk[53][5] = -11; wk[53][6] = -5; wk[53][7] = -2; wk[53][8] = 7; wk[53][9] = -9; wk[53][10] = -2; wk[53][11] = -12; wk[53][12] = 15; wk[53][13] = 9; wk[53][14] = -3; wk[53][15] = -6; 
wk[54][0] = -10; wk[54][1] = 0; wk[54][2] = -9; wk[54][3] = 3; wk[54][4] = -15; wk[54][5] = -8; wk[54][6] = 7; wk[54][7] = 2; wk[54][8] = -16; wk[54][9] = 3; wk[54][10] = -7; wk[54][11] = 11; wk[54][12] = -8; wk[54][13] = 4; wk[54][14] = 0; wk[54][15] = 15; 
wk[55][0] = -6; wk[55][1] = 0; wk[55][2] = 16; wk[55][3] = 7; wk[55][4] = 7; wk[55][5] = -9; wk[55][6] = 14; wk[55][7] = 3; wk[55][8] = 0; wk[55][9] = -1; wk[55][10] = -9; wk[55][11] = 14; wk[55][12] = -1; wk[55][13] = 7; wk[55][14] = 5; wk[55][15] = 1; 
wk[56][0] = 6; wk[56][1] = 7; wk[56][2] = 13; wk[56][3] = 9; wk[56][4] = 4; wk[56][5] = 4; wk[56][6] = -2; wk[56][7] = -11; wk[56][8] = -14; wk[56][9] = 13; wk[56][10] = -16; wk[56][11] = 3; wk[56][12] = 14; wk[56][13] = -2; wk[56][14] = -1; wk[56][15] = 0; 
wk[57][0] = -16; wk[57][1] = 6; wk[57][2] = -10; wk[57][3] = 5; wk[57][4] = 8; wk[57][5] = -13; wk[57][6] = 16; wk[57][7] = 3; wk[57][8] = 1; wk[57][9] = -3; wk[57][10] = 12; wk[57][11] = 5; wk[57][12] = -10; wk[57][13] = -14; wk[57][14] = 16; wk[57][15] = -1; 
wk[58][0] = -7; wk[58][1] = 11; wk[58][2] = 14; wk[58][3] = 6; wk[58][4] = -6; wk[58][5] = -9; wk[58][6] = 11; wk[58][7] = 5; wk[58][8] = -8; wk[58][9] = -5; wk[58][10] = 6; wk[58][11] = -8; wk[58][12] = 10; wk[58][13] = 12; wk[58][14] = 10; wk[58][15] = 1; 
wk[59][0] = -14; wk[59][1] = 12; wk[59][2] = 10; wk[59][3] = 7; wk[59][4] = -13; wk[59][5] = 1; wk[59][6] = 12; wk[59][7] = 8; wk[59][8] = 14; wk[59][9] = 10; wk[59][10] = -3; wk[59][11] = -13; wk[59][12] = -16; wk[59][13] = -3; wk[59][14] = -15; wk[59][15] = 16; 
wk[60][0] = 10; wk[60][1] = -1; wk[60][2] = 14; wk[60][3] = -6; wk[60][4] = 10; wk[60][5] = 14; wk[60][6] = 5; wk[60][7] = -8; wk[60][8] = -8; wk[60][9] = 9; wk[60][10] = 11; wk[60][11] = 8; wk[60][12] = 16; wk[60][13] = 6; wk[60][14] = -16; wk[60][15] = -12; 
wk[61][0] = -1; wk[61][1] = -11; wk[61][2] = 13; wk[61][3] = 3; wk[61][4] = -7; wk[61][5] = 15; wk[61][6] = 11; wk[61][7] = -7; wk[61][8] = -9; wk[61][9] = -10; wk[61][10] = 11; wk[61][11] = 16; wk[61][12] = -1; wk[61][13] = -5; wk[61][14] = -3; wk[61][15] = 12; 
wk[62][0] = 10; wk[62][1] = 13; wk[62][2] = -13; wk[62][3] = 13; wk[62][4] = -2; wk[62][5] = -4; wk[62][6] = -8; wk[62][7] = -3; wk[62][8] = -10; wk[62][9] = 13; wk[62][10] = -7; wk[62][11] = -8; wk[62][12] = 10; wk[62][13] = 8; wk[62][14] = 6; wk[62][15] = -1; 
wk[63][0] = -8; wk[63][1] = 11; wk[63][2] = 2; wk[63][3] = -9; wk[63][4] = -7; wk[63][5] = -14; wk[63][6] = 10; wk[63][7] = 0; wk[63][8] = 5; wk[63][9] = -16; wk[63][10] = 2; wk[63][11] = 8; wk[63][12] = 7; wk[63][13] = 13; wk[63][14] = 6; wk[63][15] = 9; 

wv[0][0] = 14; wv[0][1] = -5; wv[0][2] = 5; wv[0][3] = 8; wv[0][4] = 11; wv[0][5] = -5; wv[0][6] = 7; wv[0][7] = -13; wv[0][8] = -2; wv[0][9] = -10; wv[0][10] = 3; wv[0][11] = 11; wv[0][12] = -4; wv[0][13] = -6; wv[0][14] = 5; wv[0][15] = -5; 
wv[1][0] = 16; wv[1][1] = 9; wv[1][2] = -10; wv[1][3] = 2; wv[1][4] = 14; wv[1][5] = -16; wv[1][6] = -2; wv[1][7] = 14; wv[1][8] = -3; wv[1][9] = -12; wv[1][10] = -12; wv[1][11] = -15; wv[1][12] = -5; wv[1][13] = 4; wv[1][14] = -15; wv[1][15] = 2; 
wv[2][0] = -1; wv[2][1] = -15; wv[2][2] = -9; wv[2][3] = -5; wv[2][4] = -12; wv[2][5] = -5; wv[2][6] = -6; wv[2][7] = 13; wv[2][8] = -5; wv[2][9] = 13; wv[2][10] = -12; wv[2][11] = 0; wv[2][12] = 13; wv[2][13] = 1; wv[2][14] = -7; wv[2][15] = 2; 
wv[3][0] = 0; wv[3][1] = -7; wv[3][2] = -13; wv[3][3] = -3; wv[3][4] = 10; wv[3][5] = 7; wv[3][6] = 3; wv[3][7] = -5; wv[3][8] = 9; wv[3][9] = -5; wv[3][10] = 14; wv[3][11] = 15; wv[3][12] = 14; wv[3][13] = 15; wv[3][14] = -7; wv[3][15] = -8; 
wv[4][0] = -13; wv[4][1] = 8; wv[4][2] = -8; wv[4][3] = 7; wv[4][4] = 14; wv[4][5] = -12; wv[4][6] = 11; wv[4][7] = -8; wv[4][8] = -1; wv[4][9] = -3; wv[4][10] = 8; wv[4][11] = -7; wv[4][12] = 9; wv[4][13] = -3; wv[4][14] = -5; wv[4][15] = 8; 
wv[5][0] = 5; wv[5][1] = -7; wv[5][2] = 10; wv[5][3] = -16; wv[5][4] = 16; wv[5][5] = 2; wv[5][6] = -9; wv[5][7] = -11; wv[5][8] = -6; wv[5][9] = -11; wv[5][10] = 14; wv[5][11] = -9; wv[5][12] = -2; wv[5][13] = 12; wv[5][14] = 10; wv[5][15] = 12; 
wv[6][0] = 14; wv[6][1] = 9; wv[6][2] = -15; wv[6][3] = 13; wv[6][4] = -1; wv[6][5] = -6; wv[6][6] = -13; wv[6][7] = 3; wv[6][8] = -15; wv[6][9] = 4; wv[6][10] = -1; wv[6][11] = -7; wv[6][12] = 6; wv[6][13] = 6; wv[6][14] = -7; wv[6][15] = -7; 
wv[7][0] = 16; wv[7][1] = 6; wv[7][2] = 5; wv[7][3] = -13; wv[7][4] = 7; wv[7][5] = 14; wv[7][6] = -6; wv[7][7] = 2; wv[7][8] = 11; wv[7][9] = -6; wv[7][10] = 9; wv[7][11] = -1; wv[7][12] = 15; wv[7][13] = 15; wv[7][14] = -1; wv[7][15] = 12; 
wv[8][0] = 11; wv[8][1] = 10; wv[8][2] = 7; wv[8][3] = -4; wv[8][4] = -4; wv[8][5] = -16; wv[8][6] = 4; wv[8][7] = -5; wv[8][8] = 8; wv[8][9] = 16; wv[8][10] = -11; wv[8][11] = -10; wv[8][12] = -1; wv[8][13] = 2; wv[8][14] = 6; wv[8][15] = -16; 
wv[9][0] = 9; wv[9][1] = -8; wv[9][2] = 14; wv[9][3] = -6; wv[9][4] = 1; wv[9][5] = 12; wv[9][6] = -14; wv[9][7] = 3; wv[9][8] = -8; wv[9][9] = 6; wv[9][10] = 2; wv[9][11] = 0; wv[9][12] = 13; wv[9][13] = -6; wv[9][14] = -7; wv[9][15] = 12; 
wv[10][0] = 1; wv[10][1] = -4; wv[10][2] = -13; wv[10][3] = -13; wv[10][4] = 13; wv[10][5] = 0; wv[10][6] = 6; wv[10][7] = -1; wv[10][8] = 1; wv[10][9] = 16; wv[10][10] = 13; wv[10][11] = 5; wv[10][12] = 2; wv[10][13] = 7; wv[10][14] = -5; wv[10][15] = 11; 
wv[11][0] = -10; wv[11][1] = -11; wv[11][2] = 11; wv[11][3] = -5; wv[11][4] = 2; wv[11][5] = -4; wv[11][6] = 4; wv[11][7] = 14; wv[11][8] = -13; wv[11][9] = -15; wv[11][10] = -5; wv[11][11] = 15; wv[11][12] = -13; wv[11][13] = -7; wv[11][14] = 14; wv[11][15] = -15; 
wv[12][0] = 1; wv[12][1] = 16; wv[12][2] = -1; wv[12][3] = 7; wv[12][4] = -7; wv[12][5] = -3; wv[12][6] = -12; wv[12][7] = -13; wv[12][8] = -16; wv[12][9] = -3; wv[12][10] = 2; wv[12][11] = 8; wv[12][12] = 14; wv[12][13] = -5; wv[12][14] = 2; wv[12][15] = 2; 
wv[13][0] = -12; wv[13][1] = 11; wv[13][2] = -6; wv[13][3] = -2; wv[13][4] = -12; wv[13][5] = 10; wv[13][6] = 16; wv[13][7] = 0; wv[13][8] = -16; wv[13][9] = -12; wv[13][10] = 1; wv[13][11] = 4; wv[13][12] = 4; wv[13][13] = 6; wv[13][14] = 7; wv[13][15] = -13; 
wv[14][0] = 16; wv[14][1] = 7; wv[14][2] = -15; wv[14][3] = 6; wv[14][4] = 8; wv[14][5] = 4; wv[14][6] = 2; wv[14][7] = 6; wv[14][8] = 10; wv[14][9] = -7; wv[14][10] = 5; wv[14][11] = 11; wv[14][12] = -2; wv[14][13] = -6; wv[14][14] = 7; wv[14][15] = -5; 
wv[15][0] = -15; wv[15][1] = -12; wv[15][2] = 0; wv[15][3] = -10; wv[15][4] = 8; wv[15][5] = 4; wv[15][6] = -2; wv[15][7] = -8; wv[15][8] = 2; wv[15][9] = -13; wv[15][10] = 11; wv[15][11] = 7; wv[15][12] = 16; wv[15][13] = 15; wv[15][14] = 0; wv[15][15] = 9; 
wv[16][0] = -2; wv[16][1] = -9; wv[16][2] = 10; wv[16][3] = -14; wv[16][4] = 11; wv[16][5] = -2; wv[16][6] = 2; wv[16][7] = -15; wv[16][8] = -3; wv[16][9] = -7; wv[16][10] = 0; wv[16][11] = -8; wv[16][12] = 0; wv[16][13] = 9; wv[16][14] = 10; wv[16][15] = 4; 
wv[17][0] = -15; wv[17][1] = -6; wv[17][2] = -1; wv[17][3] = -6; wv[17][4] = -10; wv[17][5] = 7; wv[17][6] = 13; wv[17][7] = 13; wv[17][8] = 15; wv[17][9] = -5; wv[17][10] = -1; wv[17][11] = -14; wv[17][12] = -12; wv[17][13] = 14; wv[17][14] = -3; wv[17][15] = -9; 
wv[18][0] = 1; wv[18][1] = 16; wv[18][2] = -4; wv[18][3] = 3; wv[18][4] = 6; wv[18][5] = 0; wv[18][6] = 10; wv[18][7] = -12; wv[18][8] = 6; wv[18][9] = -12; wv[18][10] = -5; wv[18][11] = 5; wv[18][12] = 9; wv[18][13] = 5; wv[18][14] = -16; wv[18][15] = 3; 
wv[19][0] = -3; wv[19][1] = -16; wv[19][2] = 0; wv[19][3] = 6; wv[19][4] = 4; wv[19][5] = 10; wv[19][6] = -13; wv[19][7] = -16; wv[19][8] = 11; wv[19][9] = 11; wv[19][10] = -6; wv[19][11] = 0; wv[19][12] = 1; wv[19][13] = -1; wv[19][14] = 11; wv[19][15] = 8; 
wv[20][0] = -9; wv[20][1] = 15; wv[20][2] = -7; wv[20][3] = 14; wv[20][4] = 0; wv[20][5] = 9; wv[20][6] = 7; wv[20][7] = 14; wv[20][8] = -7; wv[20][9] = -5; wv[20][10] = -8; wv[20][11] = -11; wv[20][12] = 4; wv[20][13] = -9; wv[20][14] = -10; wv[20][15] = -11; 
wv[21][0] = 7; wv[21][1] = -11; wv[21][2] = 13; wv[21][3] = -11; wv[21][4] = 15; wv[21][5] = 9; wv[21][6] = -2; wv[21][7] = 8; wv[21][8] = -13; wv[21][9] = 15; wv[21][10] = 13; wv[21][11] = -12; wv[21][12] = -15; wv[21][13] = 11; wv[21][14] = 16; wv[21][15] = 10; 
wv[22][0] = -5; wv[22][1] = -10; wv[22][2] = -16; wv[22][3] = 4; wv[22][4] = 16; wv[22][5] = -6; wv[22][6] = 12; wv[22][7] = 8; wv[22][8] = 13; wv[22][9] = -8; wv[22][10] = 6; wv[22][11] = -16; wv[22][12] = 9; wv[22][13] = -5; wv[22][14] = -14; wv[22][15] = -6; 
wv[23][0] = 5; wv[23][1] = -9; wv[23][2] = 8; wv[23][3] = 13; wv[23][4] = 5; wv[23][5] = 5; wv[23][6] = -3; wv[23][7] = -8; wv[23][8] = 4; wv[23][9] = -8; wv[23][10] = 16; wv[23][11] = 15; wv[23][12] = -13; wv[23][13] = 10; wv[23][14] = 0; wv[23][15] = 3; 
wv[24][0] = -13; wv[24][1] = 8; wv[24][2] = -15; wv[24][3] = -11; wv[24][4] = -15; wv[24][5] = -6; wv[24][6] = 4; wv[24][7] = 14; wv[24][8] = 7; wv[24][9] = 13; wv[24][10] = -11; wv[24][11] = -4; wv[24][12] = -5; wv[24][13] = 15; wv[24][14] = 3; wv[24][15] = -13; 
wv[25][0] = -12; wv[25][1] = -9; wv[25][2] = -1; wv[25][3] = -12; wv[25][4] = 4; wv[25][5] = 2; wv[25][6] = -12; wv[25][7] = 3; wv[25][8] = 3; wv[25][9] = -3; wv[25][10] = -16; wv[25][11] = 1; wv[25][12] = -11; wv[25][13] = 10; wv[25][14] = -14; wv[25][15] = -10; 
wv[26][0] = 14; wv[26][1] = 10; wv[26][2] = -5; wv[26][3] = -6; wv[26][4] = -10; wv[26][5] = 3; wv[26][6] = -2; wv[26][7] = -12; wv[26][8] = 16; wv[26][9] = 15; wv[26][10] = -1; wv[26][11] = 6; wv[26][12] = 16; wv[26][13] = 13; wv[26][14] = 13; wv[26][15] = -10; 
wv[27][0] = 11; wv[27][1] = 12; wv[27][2] = -1; wv[27][3] = -1; wv[27][4] = 10; wv[27][5] = 6; wv[27][6] = 3; wv[27][7] = -11; wv[27][8] = 14; wv[27][9] = -6; wv[27][10] = 1; wv[27][11] = 13; wv[27][12] = 1; wv[27][13] = -16; wv[27][14] = 13; wv[27][15] = 1; 
wv[28][0] = 9; wv[28][1] = -13; wv[28][2] = 0; wv[28][3] = 2; wv[28][4] = 12; wv[28][5] = 5; wv[28][6] = 7; wv[28][7] = 8; wv[28][8] = -4; wv[28][9] = -7; wv[28][10] = 4; wv[28][11] = 6; wv[28][12] = -14; wv[28][13] = 1; wv[28][14] = -11; wv[28][15] = 10; 
wv[29][0] = 5; wv[29][1] = 3; wv[29][2] = 11; wv[29][3] = -11; wv[29][4] = -5; wv[29][5] = 12; wv[29][6] = 16; wv[29][7] = 2; wv[29][8] = 14; wv[29][9] = 1; wv[29][10] = 2; wv[29][11] = -14; wv[29][12] = 1; wv[29][13] = -11; wv[29][14] = 10; wv[29][15] = -8; 
wv[30][0] = -2; wv[30][1] = -10; wv[30][2] = 2; wv[30][3] = 1; wv[30][4] = 2; wv[30][5] = -12; wv[30][6] = -6; wv[30][7] = -3; wv[30][8] = 9; wv[30][9] = -9; wv[30][10] = 7; wv[30][11] = 16; wv[30][12] = -5; wv[30][13] = 2; wv[30][14] = -10; wv[30][15] = 7; 
wv[31][0] = 7; wv[31][1] = 4; wv[31][2] = 11; wv[31][3] = -10; wv[31][4] = 11; wv[31][5] = 1; wv[31][6] = 5; wv[31][7] = 10; wv[31][8] = -3; wv[31][9] = -7; wv[31][10] = -11; wv[31][11] = 13; wv[31][12] = -8; wv[31][13] = -1; wv[31][14] = 7; wv[31][15] = -12; 
wv[32][0] = -9; wv[32][1] = -1; wv[32][2] = -15; wv[32][3] = 3; wv[32][4] = -12; wv[32][5] = 9; wv[32][6] = 2; wv[32][7] = -11; wv[32][8] = -14; wv[32][9] = -13; wv[32][10] = 15; wv[32][11] = 9; wv[32][12] = 3; wv[32][13] = 15; wv[32][14] = 9; wv[32][15] = 16; 
wv[33][0] = 15; wv[33][1] = 13; wv[33][2] = 0; wv[33][3] = 7; wv[33][4] = -2; wv[33][5] = 10; wv[33][6] = -6; wv[33][7] = -2; wv[33][8] = -1; wv[33][9] = 13; wv[33][10] = 16; wv[33][11] = -5; wv[33][12] = 15; wv[33][13] = 1; wv[33][14] = 3; wv[33][15] = -9; 
wv[34][0] = -3; wv[34][1] = 16; wv[34][2] = 9; wv[34][3] = 4; wv[34][4] = 7; wv[34][5] = -16; wv[34][6] = -14; wv[34][7] = 15; wv[34][8] = -15; wv[34][9] = -2; wv[34][10] = -3; wv[34][11] = -16; wv[34][12] = 13; wv[34][13] = -4; wv[34][14] = -5; wv[34][15] = 3; 
wv[35][0] = -1; wv[35][1] = -16; wv[35][2] = 15; wv[35][3] = 1; wv[35][4] = -3; wv[35][5] = 6; wv[35][6] = 8; wv[35][7] = -4; wv[35][8] = -8; wv[35][9] = 5; wv[35][10] = -16; wv[35][11] = 10; wv[35][12] = -13; wv[35][13] = 5; wv[35][14] = 11; wv[35][15] = -16; 
wv[36][0] = -6; wv[36][1] = -3; wv[36][2] = 11; wv[36][3] = -12; wv[36][4] = 7; wv[36][5] = 13; wv[36][6] = -5; wv[36][7] = 9; wv[36][8] = -6; wv[36][9] = -10; wv[36][10] = 16; wv[36][11] = -1; wv[36][12] = -11; wv[36][13] = 10; wv[36][14] = 14; wv[36][15] = 7; 
wv[37][0] = 12; wv[37][1] = 0; wv[37][2] = -7; wv[37][3] = -14; wv[37][4] = 1; wv[37][5] = -8; wv[37][6] = 3; wv[37][7] = 5; wv[37][8] = -3; wv[37][9] = -1; wv[37][10] = 13; wv[37][11] = 5; wv[37][12] = -5; wv[37][13] = -10; wv[37][14] = 1; wv[37][15] = -9; 
wv[38][0] = 15; wv[38][1] = 8; wv[38][2] = 8; wv[38][3] = -1; wv[38][4] = 1; wv[38][5] = -4; wv[38][6] = -5; wv[38][7] = 4; wv[38][8] = -2; wv[38][9] = 9; wv[38][10] = -1; wv[38][11] = -16; wv[38][12] = 7; wv[38][13] = 12; wv[38][14] = 6; wv[38][15] = 3; 
wv[39][0] = -14; wv[39][1] = 0; wv[39][2] = -5; wv[39][3] = 14; wv[39][4] = 15; wv[39][5] = 8; wv[39][6] = -6; wv[39][7] = 0; wv[39][8] = 11; wv[39][9] = -12; wv[39][10] = 11; wv[39][11] = -13; wv[39][12] = -15; wv[39][13] = -16; wv[39][14] = 5; wv[39][15] = -8; 
wv[40][0] = 8; wv[40][1] = -5; wv[40][2] = 14; wv[40][3] = 10; wv[40][4] = -15; wv[40][5] = 3; wv[40][6] = -6; wv[40][7] = 5; wv[40][8] = 15; wv[40][9] = -16; wv[40][10] = 1; wv[40][11] = 6; wv[40][12] = 10; wv[40][13] = -4; wv[40][14] = -6; wv[40][15] = -16; 
wv[41][0] = 1; wv[41][1] = -7; wv[41][2] = -6; wv[41][3] = 9; wv[41][4] = -1; wv[41][5] = -16; wv[41][6] = -1; wv[41][7] = -7; wv[41][8] = -10; wv[41][9] = 6; wv[41][10] = -12; wv[41][11] = 7; wv[41][12] = -6; wv[41][13] = 3; wv[41][14] = -2; wv[41][15] = -15; 
wv[42][0] = -3; wv[42][1] = 5; wv[42][2] = -2; wv[42][3] = -11; wv[42][4] = -13; wv[42][5] = 7; wv[42][6] = 5; wv[42][7] = -7; wv[42][8] = -5; wv[42][9] = -7; wv[42][10] = -13; wv[42][11] = -13; wv[42][12] = -9; wv[42][13] = -11; wv[42][14] = -6; wv[42][15] = -3; 
wv[43][0] = -1; wv[43][1] = 11; wv[43][2] = 7; wv[43][3] = 5; wv[43][4] = 0; wv[43][5] = -1; wv[43][6] = 3; wv[43][7] = -8; wv[43][8] = -7; wv[43][9] = -14; wv[43][10] = 15; wv[43][11] = 4; wv[43][12] = -15; wv[43][13] = 11; wv[43][14] = 15; wv[43][15] = -4; 
wv[44][0] = 13; wv[44][1] = 10; wv[44][2] = 8; wv[44][3] = -14; wv[44][4] = -10; wv[44][5] = -5; wv[44][6] = -2; wv[44][7] = 14; wv[44][8] = 14; wv[44][9] = 14; wv[44][10] = -14; wv[44][11] = -4; wv[44][12] = -16; wv[44][13] = -2; wv[44][14] = -10; wv[44][15] = -14; 
wv[45][0] = 3; wv[45][1] = 3; wv[45][2] = -2; wv[45][3] = 10; wv[45][4] = -11; wv[45][5] = -15; wv[45][6] = 11; wv[45][7] = 4; wv[45][8] = -14; wv[45][9] = 6; wv[45][10] = 1; wv[45][11] = -4; wv[45][12] = 4; wv[45][13] = 16; wv[45][14] = 12; wv[45][15] = 8; 
wv[46][0] = 16; wv[46][1] = 3; wv[46][2] = 1; wv[46][3] = 11; wv[46][4] = 1; wv[46][5] = 3; wv[46][6] = 15; wv[46][7] = -5; wv[46][8] = 10; wv[46][9] = 15; wv[46][10] = -3; wv[46][11] = 16; wv[46][12] = -15; wv[46][13] = -2; wv[46][14] = -4; wv[46][15] = 2; 
wv[47][0] = 15; wv[47][1] = 6; wv[47][2] = -10; wv[47][3] = -7; wv[47][4] = 15; wv[47][5] = 6; wv[47][6] = -4; wv[47][7] = -6; wv[47][8] = 7; wv[47][9] = 14; wv[47][10] = 16; wv[47][11] = 3; wv[47][12] = 0; wv[47][13] = -13; wv[47][14] = -7; wv[47][15] = -15; 
wv[48][0] = -10; wv[48][1] = -13; wv[48][2] = 0; wv[48][3] = -8; wv[48][4] = -11; wv[48][5] = 15; wv[48][6] = 5; wv[48][7] = -4; wv[48][8] = 12; wv[48][9] = -4; wv[48][10] = -7; wv[48][11] = -4; wv[48][12] = -3; wv[48][13] = 5; wv[48][14] = 5; wv[48][15] = -8; 
wv[49][0] = -14; wv[49][1] = -6; wv[49][2] = 5; wv[49][3] = 8; wv[49][4] = -1; wv[49][5] = -14; wv[49][6] = 5; wv[49][7] = -6; wv[49][8] = -16; wv[49][9] = 2; wv[49][10] = -8; wv[49][11] = -1; wv[49][12] = -13; wv[49][13] = 4; wv[49][14] = 5; wv[49][15] = 13; 
wv[50][0] = 2; wv[50][1] = 16; wv[50][2] = 9; wv[50][3] = 13; wv[50][4] = -9; wv[50][5] = -8; wv[50][6] = -11; wv[50][7] = 14; wv[50][8] = -5; wv[50][9] = -11; wv[50][10] = -7; wv[50][11] = -12; wv[50][12] = -9; wv[50][13] = -11; wv[50][14] = -8; wv[50][15] = -6; 
wv[51][0] = -14; wv[51][1] = -13; wv[51][2] = -2; wv[51][3] = -3; wv[51][4] = -1; wv[51][5] = -13; wv[51][6] = -10; wv[51][7] = 8; wv[51][8] = 16; wv[51][9] = -9; wv[51][10] = -8; wv[51][11] = 3; wv[51][12] = -3; wv[51][13] = -16; wv[51][14] = -3; wv[51][15] = 12; 
wv[52][0] = -4; wv[52][1] = -9; wv[52][2] = 14; wv[52][3] = 3; wv[52][4] = 11; wv[52][5] = 6; wv[52][6] = 15; wv[52][7] = -10; wv[52][8] = 6; wv[52][9] = -12; wv[52][10] = -15; wv[52][11] = 7; wv[52][12] = 8; wv[52][13] = 4; wv[52][14] = -14; wv[52][15] = -2; 
wv[53][0] = 11; wv[53][1] = 2; wv[53][2] = -15; wv[53][3] = -15; wv[53][4] = 7; wv[53][5] = 5; wv[53][6] = -11; wv[53][7] = 2; wv[53][8] = -16; wv[53][9] = 0; wv[53][10] = 2; wv[53][11] = -2; wv[53][12] = 11; wv[53][13] = 4; wv[53][14] = 3; wv[53][15] = -7; 
wv[54][0] = 13; wv[54][1] = -2; wv[54][2] = 13; wv[54][3] = -4; wv[54][4] = -13; wv[54][5] = 13; wv[54][6] = -9; wv[54][7] = 10; wv[54][8] = 2; wv[54][9] = 0; wv[54][10] = 15; wv[54][11] = 3; wv[54][12] = 13; wv[54][13] = 6; wv[54][14] = 0; wv[54][15] = 14; 
wv[55][0] = 2; wv[55][1] = -11; wv[55][2] = 3; wv[55][3] = 10; wv[55][4] = 0; wv[55][5] = 7; wv[55][6] = 12; wv[55][7] = 2; wv[55][8] = -11; wv[55][9] = -3; wv[55][10] = -13; wv[55][11] = 14; wv[55][12] = 5; wv[55][13] = -11; wv[55][14] = 3; wv[55][15] = -12; 
wv[56][0] = -3; wv[56][1] = -2; wv[56][2] = -13; wv[56][3] = -14; wv[56][4] = -13; wv[56][5] = -11; wv[56][6] = 10; wv[56][7] = 2; wv[56][8] = 11; wv[56][9] = -2; wv[56][10] = -3; wv[56][11] = 13; wv[56][12] = 0; wv[56][13] = 14; wv[56][14] = 12; wv[56][15] = 14; 
wv[57][0] = 2; wv[57][1] = 9; wv[57][2] = 4; wv[57][3] = 14; wv[57][4] = -5; wv[57][5] = 5; wv[57][6] = 6; wv[57][7] = -13; wv[57][8] = 2; wv[57][9] = -8; wv[57][10] = 13; wv[57][11] = -13; wv[57][12] = 12; wv[57][13] = -8; wv[57][14] = 1; wv[57][15] = -10; 
wv[58][0] = -2; wv[58][1] = 10; wv[58][2] = -16; wv[58][3] = 16; wv[58][4] = 8; wv[58][5] = -11; wv[58][6] = -10; wv[58][7] = 4; wv[58][8] = -15; wv[58][9] = -7; wv[58][10] = -13; wv[58][11] = -9; wv[58][12] = -3; wv[58][13] = -5; wv[58][14] = 1; wv[58][15] = -9; 
wv[59][0] = -13; wv[59][1] = 3; wv[59][2] = 1; wv[59][3] = -14; wv[59][4] = -15; wv[59][5] = 4; wv[59][6] = 8; wv[59][7] = 4; wv[59][8] = -5; wv[59][9] = -11; wv[59][10] = 1; wv[59][11] = 8; wv[59][12] = 8; wv[59][13] = -1; wv[59][14] = -11; wv[59][15] = 14; 
wv[60][0] = 8; wv[60][1] = 15; wv[60][2] = 1; wv[60][3] = -13; wv[60][4] = 5; wv[60][5] = 11; wv[60][6] = 0; wv[60][7] = 4; wv[60][8] = 14; wv[60][9] = -16; wv[60][10] = -15; wv[60][11] = 0; wv[60][12] = 3; wv[60][13] = 8; wv[60][14] = 11; wv[60][15] = -4; 
wv[61][0] = -6; wv[61][1] = 12; wv[61][2] = -14; wv[61][3] = -9; wv[61][4] = 6; wv[61][5] = -14; wv[61][6] = 4; wv[61][7] = 3; wv[61][8] = 6; wv[61][9] = -5; wv[61][10] = -2; wv[61][11] = 15; wv[61][12] = -10; wv[61][13] = 1; wv[61][14] = 6; wv[61][15] = -12; 
wv[62][0] = 15; wv[62][1] = -7; wv[62][2] = 16; wv[62][3] = 2; wv[62][4] = 4; wv[62][5] = 10; wv[62][6] = 4; wv[62][7] = -9; wv[62][8] = 7; wv[62][9] = -2; wv[62][10] = -11; wv[62][11] = 4; wv[62][12] = -2; wv[62][13] = 15; wv[62][14] = 2; wv[62][15] = 14; 
wv[63][0] = -3; wv[63][1] = 1; wv[63][2] = -12; wv[63][3] = -4; wv[63][4] = 4; wv[63][5] = -9; wv[63][6] = -1; wv[63][7] = 4; wv[63][8] = -4; wv[63][9] = -15; wv[63][10] = 2; wv[63][11] = 7; wv[63][12] = 8; wv[63][13] = 2; wv[63][14] = 8; wv[63][15] = -6; 


    //Iteratively interfacing 64 elements of the weight column across three interfaces - 16 times
    rule load_weights (start1 == 0);
        if (stepq < (fromInteger(w_cols)+1)) 
        begin
            dut.get_weightsq(wq[0][stepq], wq[1][stepq], wq[2][stepq], wq[3][stepq], wq[4][stepq], wq[5][stepq], wq[6][stepq], wq[7][stepq], wq[8][stepq], wq[9][stepq], wq[10][stepq], wq[11][stepq], wq[12][stepq], wq[13][stepq], wq[14][stepq], wq[15][stepq], wq[16][stepq], wq[17][stepq], wq[18][stepq], wq[19][stepq], wq[20][stepq], wq[21][stepq], wq[22][stepq], wq[23][stepq], wq[24][stepq], wq[25][stepq], wq[26][stepq], wq[27][stepq], wq[28][stepq], wq[29][stepq], wq[30][stepq], wq[31][stepq], wq[32][stepq], wq[33][stepq], wq[34][stepq], wq[35][stepq], wq[36][stepq], wq[37][stepq], wq[38][stepq], wq[39][stepq], wq[40][stepq], wq[41][stepq], wq[42][stepq], wq[43][stepq], wq[44][stepq], wq[45][stepq], wq[46][stepq], wq[47][stepq], wq[48][stepq], wq[49][stepq], wq[50][stepq], wq[51][stepq], wq[52][stepq], wq[53][stepq], wq[54][stepq], wq[55][stepq], wq[56][stepq], wq[57][stepq], wq[58][stepq], wq[59][stepq], wq[60][stepq], wq[61][stepq], wq[62][stepq], wq[63][stepq]);
            dut.get_weightsk(wk[0][stepq], wk[1][stepq], wk[2][stepq], wk[3][stepq], wk[4][stepq], wk[5][stepq], wk[6][stepq], wk[7][stepq], wk[8][stepq], wk[9][stepq], wk[10][stepq], wk[11][stepq], wk[12][stepq], wk[13][stepq], wk[14][stepq], wk[15][stepq], wk[16][stepq], wk[17][stepq], wk[18][stepq], wk[19][stepq], wk[20][stepq], wk[21][stepq], wk[22][stepq], wk[23][stepq], wk[24][stepq], wk[25][stepq], wk[26][stepq], wk[27][stepq], wk[28][stepq], wk[29][stepq], wk[30][stepq], wk[31][stepq], wk[32][stepq], wk[33][stepq], wk[34][stepq], wk[35][stepq], wk[36][stepq], wk[37][stepq], wk[38][stepq], wk[39][stepq], wk[40][stepq], wk[41][stepq], wk[42][stepq], wk[43][stepq], wk[44][stepq], wk[45][stepq], wk[46][stepq], wk[47][stepq], wk[48][stepq], wk[49][stepq], wk[50][stepq], wk[51][stepq], wk[52][stepq], wk[53][stepq], wk[54][stepq], wk[55][stepq], wk[56][stepq], wk[57][stepq], wk[58][stepq], wk[59][stepq], wk[60][stepq], wk[61][stepq], wk[62][stepq], wk[63][stepq]);
            dut.get_weightsv(wv[0][stepq], wv[1][stepq], wv[2][stepq], wv[3][stepq], wv[4][stepq], wv[5][stepq], wv[6][stepq], wv[7][stepq], wv[8][stepq], wv[9][stepq], wv[10][stepq], wv[11][stepq], wv[12][stepq], wv[13][stepq], wv[14][stepq], wv[15][stepq], wv[16][stepq], wv[17][stepq], wv[18][stepq], wv[19][stepq], wv[20][stepq], wv[21][stepq], wv[22][stepq], wv[23][stepq], wv[24][stepq], wv[25][stepq], wv[26][stepq], wv[27][stepq], wv[28][stepq], wv[29][stepq], wv[30][stepq], wv[31][stepq], wv[32][stepq], wv[33][stepq], wv[34][stepq], wv[35][stepq], wv[36][stepq], wv[37][stepq], wv[38][stepq], wv[39][stepq], wv[40][stepq], wv[41][stepq], wv[42][stepq], wv[43][stepq], wv[44][stepq], wv[45][stepq], wv[46][stepq], wv[47][stepq], wv[48][stepq], wv[49][stepq], wv[50][stepq], wv[51][stepq], wv[52][stepq], wv[53][stepq], wv[54][stepq], wv[55][stepq], wv[56][stepq], wv[57][stepq], wv[58][stepq], wv[59][stepq], wv[60][stepq], wv[61][stepq], wv[62][stepq], wv[63][stepq]);
            start1 <= 0;
            stepq <= stepq + 1;
        end
        else 
            begin
            start1 <= 2;
        end
    endrule
        

    //Iteratively interfacing 64 elements of the Input rows - 16 times
    rule load_inputs (start1 == 2);
    if(stepx < fromInteger(in_rows))
    begin
        dut.get_inputs(x[stepx][0], x[stepx][1], x[stepx][2], x[stepx][3], x[stepx][4], x[stepx][5], x[stepx][6], x[stepx][7], x[stepx][8], x[stepx][9], x[stepx][10], x[stepx][11], x[stepx][12], x[stepx][13], x[stepx][14], x[stepx][15], x[stepx][16], x[stepx][17], x[stepx][18], x[stepx][19], x[stepx][20], x[stepx][21], x[stepx][22], x[stepx][23], x[stepx][24], x[stepx][25], x[stepx][26], x[stepx][27], x[stepx][28], x[stepx][29], x[stepx][30], x[stepx][31], x[stepx][32], x[stepx][33], x[stepx][34], x[stepx][35], x[stepx][36], x[stepx][37], x[stepx][38], x[stepx][39], x[stepx][40], x[stepx][41], x[stepx][42], x[stepx][43], x[stepx][44], x[stepx][45], x[stepx][46], x[stepx][47], x[stepx][48], x[stepx][49], x[stepx][50], x[stepx][51], x[stepx][52], x[stepx][53], x[stepx][54], x[stepx][55], x[stepx][56], x[stepx][57], x[stepx][58], x[stepx][59], x[stepx][60], x[stepx][61], x[stepx][62], x[stepx][63]); 
        start1 <= 2;
        stepx <= stepx + 1;
    end
    else 
        start1 <= 3;
    endrule

    //To capture the completion of the computation
    rule get_output (start1 == 3);
        let done = dut.get_output();
        $display("output: %b",done);
        $finish(0);
    endrule

endmodule
endpackage
